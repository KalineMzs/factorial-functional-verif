package yarvi_tb_cfg_pkg;
    parameter IN_DATA_WD = 4;
    parameter OUT_DATA_WD = 46;
endpackage
