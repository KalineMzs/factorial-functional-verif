package factorial_tb_cfg_pkg;
    parameter IN_DATA_WD = 32;
    parameter OUT_DATA_WD = 32;
endpackage
