package factorial_tb_cfg_pkg;
    parameter IN_DATA_WD = 3;
    parameter OUT_DATA_WD = 16;
endpackage
